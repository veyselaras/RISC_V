LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_PROGRAM_COUNTER IS
END TB_PROGRAM_COUNTER;

ARCHITECTURE TEST OF TB_PROGRAM_COUNTER IS


	-- CLOCK PERIYODU (10 NS = 100 MHZ CLOCK)
	
	SIGNAL CLK_TB		: STD_LOGIC := '0';
	SIGNAL RST_TB		: STD_LOGIC := '0';
	SIGNAL PC_IN_TB		: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL PC_OUT_TB	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	CONSTANT CLK_PERIOD : TIME := 10 NS;

BEGIN
	
	CLK_PROCESS:PROCESS
	BEGIN
		WHILE NOW < 100 NS LOOP  -- 100 NS SIMÜLASYON SÜRESI
            CLK_TB <= '0';
            WAIT FOR CLK_PERIOD / 2;  -- YARı PERIYOT
            CLK_TB <= '1';
            WAIT FOR CLK_PERIOD / 2;
        END LOOP;
        WAIT;
	END PROCESS;
	
	TB_PROCESS:PROCESS
	BEGIN 

		RST_TB		<= '0';
		WAIT FOR CLK_PERIOD;
		
		RST_TB		<= '1';
		WAIT FOR CLK_PERIOD;
		
		PC_IN_TB		<= X"11110000";
		WAIT FOR CLK_PERIOD;
		
		PC_IN_TB		<= X"AABB0101";
		WAIT FOR CLK_PERIOD;
		
		PC_IN_TB		<= X"CCCC0101";
		WAIT FOR CLK_PERIOD;

		PC_IN_TB		<= X"00000101";
		WAIT FOR CLK_PERIOD;
		
		RST_TB 		<= '0';
      WAIT FOR CLK_PERIOD;
		
      RST_TB		<= '1';
      WAIT FOR CLK_PERIOD;
		
		PC_IN_TB		<= X"12345678";
      WAIT FOR CLK_PERIOD;
		
		WAIT;
	END PROCESS;
	
	UUT: ENTITY WORK.PROGRAM_COUNTER
	PORT MAP (
		CLK		=> CLK_TB,
		RST		=> RST_TB,
		PC_IN		=> PC_IN_TB,
		PC_OUT	=> PC_OUT_TB
	);
	
END TEST;