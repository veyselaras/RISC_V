LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_REGISTER_FILE IS
END TB_REGISTER_FILE;

ARCHITECTURE TEST OF TB_REGISTER_FILE IS 

	SIGNAL TB_CLK					: STD_LOGIC := '0';
	
	SIGNAL TB_READ_REGISTER_1	: STD_LOGIC_VECTOR(4 DOWNTO 0) := (others => '0');
	SIGNAL TB_READ_REGISTER_2	: STD_LOGIC_VECTOR(4 DOWNTO 0) := (others => '0');
	SIGNAL TB_WRITE_REGISTER	: STD_LOGIC_VECTOR(4 DOWNTO 0) := (others => '0');
	SIGNAL TB_WRITE_DATA			: STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
	
	SIGNAL TB_CONTROL_WRITE		: STD_LOGIC := '0';
	
	SIGNAL TB_O_READ_DATA_1		: STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
	SIGNAL TB_O_READ_DATA_2		: STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
	
	CONSTANT CLK_PERIOD			 : TIME := 10 NS;
	
BEGIN
	UUT: ENTITY WORK.REGISTER_FILE
	PORT MAP
	(
		CLK					=> TB_CLK,
	
        I_READ_REGISTER_1	=> TB_READ_REGISTER_1,
        I_READ_REGISTER_2   => TB_READ_REGISTER_2,
        I_WRITE_REGISTER    => TB_WRITE_REGISTER,
        I_WRITE_DATA        => TB_WRITE_DATA,
		
        I_CONTROL_WRITE     => TB_CONTROL_WRITE,

        O_READ_DATA_1       => TB_O_READ_DATA_1,
        O_READ_DATA_2       => TB_O_READ_DATA_2
	);
	
	CLK_GEN: PROCESS
    BEGIN
        WHILE NOW<140NS LOOP
            TB_CLK <= '0';                    -- SAAT SINYALI DÜŞÜK
            WAIT FOR CLK_PERIOD/2;            -- YARıM PERIYOT BEKLEME
            TB_CLK <= '1';                    -- SAAT SINYALI YÜKSEK
            WAIT FOR CLK_PERIOD/2;            -- YARıM PERIYOT BEKLEME
        END LOOP;
    END PROCESS CLK_GEN;
	
	TEST_PROCESS: PROCESS
	BEGIN
		TB_READ_REGISTER_1	<= "00100";
		TB_READ_REGISTER_2	<= "00001";
		TB_WRITE_REGISTER	<= "11111";
		TB_WRITE_DATA		<= X"0000FFFF";
		
		TB_CONTROL_WRITE	<= '0';
		
		WAIT FOR CLK_PERIOD*2;
		
		TB_READ_REGISTER_1	<= "00000";
		TB_READ_REGISTER_2	<= "01001";
		TB_WRITE_REGISTER	<= "10111";
		TB_WRITE_DATA		<= X"0000FFFF";
		
		TB_CONTROL_WRITE	<= '1';
		
		WAIT FOR CLK_PERIOD*2;
		
		
		TB_READ_REGISTER_1	<= "00010";
		TB_READ_REGISTER_2	<= "10000";
		TB_WRITE_REGISTER	<= "11110";
		TB_WRITE_DATA		<= X"0000FFFF";
		
		TB_CONTROL_WRITE	<= '0';
		
		WAIT FOR CLK_PERIOD*2;
		
		
		TB_READ_REGISTER_1	<= "00100";
		TB_READ_REGISTER_2	<= "00001";
		TB_WRITE_REGISTER	<= "11110";
		TB_WRITE_DATA		<= X"0000FFFC";
		
		TB_CONTROL_WRITE	<= '1';
		
		WAIT FOR CLK_PERIOD*2;
		
		TB_READ_REGISTER_1	<= "01000";
		TB_READ_REGISTER_2	<= "01001";
		TB_WRITE_REGISTER	<= "11111";
		TB_WRITE_DATA		<= X"0000FAAF";
		
		TB_CONTROL_WRITE	<= '0';
		
		WAIT FOR CLK_PERIOD*2;
		
		TB_READ_REGISTER_1	<= "01000";
		TB_READ_REGISTER_2	<= "01001";
		TB_WRITE_REGISTER	<= "10001";
		TB_WRITE_DATA		<= X"0000FAAF";
		
		TB_CONTROL_WRITE	<= '1';
		
		WAIT FOR CLK_PERIOD*2;
		
		TB_READ_REGISTER_1	<= "11100";
		TB_READ_REGISTER_2	<= "11001";
		TB_WRITE_REGISTER	<= "11111";
		TB_WRITE_DATA		<= X"FFFFFFFF";
		
		TB_CONTROL_WRITE	<= '0';
		
		WAIT FOR CLK_PERIOD*2;
		
		WAIT;
	END PROCESS TEST_PROCESS;
	
END TEST;