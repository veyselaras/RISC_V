LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_INSTRUCTION_MEMORY IS
END TB_INSTRUCTION_MEMORY;

ARCHITECTURE TEST OF TB_INSTRUCTION_MEMORY IS

SIGNAL CLK_TB			: STD_LOGIC;
SIGNAL I_ADDRESS_TB		: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL O_INSTRUCTION_TB	: STD_LOGIC_VECTOR(31 DOWNTO 0);

constant CLK_PERIOD : time := 10 ns;

BEGIN
	
CLK_PROCESS:PROCESS
	BEGIN
		WHILE NOW < 100 NS LOOP  -- 100 NS SIMÜLASYON SÜRESI
            CLK_TB <= '0';
            WAIT FOR CLK_PERIOD / 2;  -- YARı PERIYOT
            CLK_TB <= '1';
            WAIT FOR CLK_PERIOD / 2;
        END LOOP;
        WAIT;
	END PROCESS;
	
TB_PROCESS:PROCESS
BEGIN
	
	I_ADDRESS_TB	<= X"00000000";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000004";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000008";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"0000000C";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000010";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000004";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000010";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"0000000C";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000010";
	WAIT FOR CLK_PERIOD;
	
	I_ADDRESS_TB	<= X"00000008";
	WAIT FOR CLK_PERIOD;
	
	WAIT;
END PROCESS;
	
	UUT: ENTITY WORK.INSTRUCTION_MEMORY
	PORT MAP (
		CLK				=> CLK_TB,
		I_ADDRESS		=> I_ADDRESS_TB,
		O_INSTRUCTION	=> O_INSTRUCTION_TB
	);
	
END TEST;